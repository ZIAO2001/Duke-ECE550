module connector(in0,out1);
	input [31:0] in0;
	output [31:0] out1;
	assign out1 = in0;
endmodule
